library verilog;
use verilog.vl_types.all;
entity ALU_4BIT_TB is
end ALU_4BIT_TB;
