library verilog;
use verilog.vl_types.all;
entity DEMO_TB_RIP is
end DEMO_TB_RIP;
