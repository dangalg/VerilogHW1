library verilog;
use verilog.vl_types.all;
entity DEMO_TB is
end DEMO_TB;
