library verilog;
use verilog.vl_types.all;
entity ALU_1BIT_TB is
end ALU_1BIT_TB;
