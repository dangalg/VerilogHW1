library verilog;
use verilog.vl_types.all;
entity DEMO_TB_FAS is
end DEMO_TB_FAS;
