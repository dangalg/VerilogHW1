library verilog;
use verilog.vl_types.all;
entity RIP_FAS_TB is
end RIP_FAS_TB;
