library verilog;
use verilog.vl_types.all;
entity FULLADDERTB is
    generic(
        delay           : integer := 15
    );
end FULLADDERTB;
