// Code your testbench here
// or browse Examples

`include "mux4_tb.sv"
`include "rip_fas_tb.sv"
`include "alu_4bit_tb.sv"
