module alu_1bit(s, cout, a, b, cin, s_op);
  input a, b, cin, s_op;
  output cout, s;
  parameter Tpd = 1;
    mux4on1
endmodule
