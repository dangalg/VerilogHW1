library verilog;
use verilog.vl_types.all;
entity MUX4_TB is
end MUX4_TB;
